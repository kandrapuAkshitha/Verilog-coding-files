module tb_down_con;
reg clk,rst;
wire [3:0] count;

down_con s(clk,rst,count);

initial clk=0;
always #5 clk =~clk;

initial begin
   rst=1;
  #10;rst=0;
   $monitor (clk,rst,count);
    #250;
   $stop;
  end
endmodule
