module complement_1s(
input [3:0] a,
output [3:0] comp);

assign comp=~a;
endmodule

