module Msb_prio_enc(
input [3:0] in,
output reg[1:0] y);

always @(*) begin
 casez(in)
  4'b1??? : y=2'b11;
  4'b01?? : y=2'b10;
  4'b001? : y=2'b01;
  4'b0001 : y=2'b00;
   default :y=2'bxx;
 endcase
 end
endmodule

